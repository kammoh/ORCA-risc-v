../../wishbone/wb_arbiter.vhd