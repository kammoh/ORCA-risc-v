library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity execute is
  generic(
	 REGISTER_SIZE			: positive;
	 REGISTER_NAME_SIZE	: positive;
	 INSTRUCTION_SIZE		: positive;
	 SIGN_EXTENSION_SIZE : positive);
  port(
	 clk	 : in std_logic;
	 reset : in std_logic;

	 pc_next		 : in std_logic_vector(REGISTER_SIZE-1 downto 0);
	 pc_current	 : in std_logic_vector(REGISTER_SIZE-1 downto 0);
	 instruction : in std_logic_vector(INSTRUCTION_SIZE-1 downto 0);

	 rs1_data		 : in std_logic_vector(REGISTER_SIZE-1 downto 0);
	 rs2_data		 : in std_logic_vector(REGISTER_SIZE-1 downto 0);
	 sign_extension : in std_logic_vector(SIGN_EXTENSION_SIZE-1 downto 0);

	 wb_sel	: inout std_logic_vector(REGISTER_NAME_SIZE-1 downto 0);
	 wb_data : inout std_logic_vector(REGISTER_SIZE-1 downto 0);
	 wb_en	: inout std_logic;

	 predict_corr	  : out std_logic_vector(REGISTER_SIZE-1 downto 0);
	 predict_corr_en : out std_logic);
end;

architecture behavioural of execute is

  alias rd : std_logic_vector(REGISTER_NAME_SIZE-1 downto 0) is
	 instruction(11 downto 7);
  alias rs1 : std_logic_vector(REGISTER_NAME_SIZE-1 downto 0) is
	 instruction(19 downto 15);
  alias rs2 : std_logic_vector(REGISTER_NAME_SIZE-1 downto 0) is
	 instruction(24 downto 20);





  -- various writeback sources
  signal br_data_out	 : std_logic_vector(REGISTER_SIZE-1 downto 0);
  signal alu_data_out : std_logic_vector(REGISTER_SIZE-1 downto 0);
  signal ld_data_out	 : std_logic_vector(REGISTER_SIZE-1 downto 0);
  signal br_data_en	 : std_logic;
  signal alu_data_en	 : std_logic;
  signal ld_data_en	 : std_logic;

  signal writeback_1hot : std_logic_vector(2 downto 0);

  signal bad_predict : std_logic;
  signal new_pc		: std_logic_vector(REGISTER_SIZE-1 downto 0);


  component arithmetic_unit is
	 generic (
		INSTRUCTION_SIZE	  : integer;
		REGISTER_SIZE		  : integer;
		SIGN_EXTENSION_SIZE : integer);
	 port (
		clk				: in	std_logic;
		rs1_data			: in	std_logic_vector(REGISTER_SIZE-1 downto 0);
		rs2_data			: in	std_logic_vector(REGISTER_SIZE-1 downto 0);
		instruction		: in	std_logic_vector(INSTRUCTION_SIZE-1 downto 0);
		sign_extension : in	std_logic_vector(SIGN_EXTENSION_SIZE-1 downto 0);
		data_out			: out std_logic_vector(REGISTER_SIZE-1 downto 0);
		data_enable		: out std_logic);
  end component arithmetic_unit;

  component branch_unit is
	 generic (
		REGISTER_SIZE		  : integer;
		INSTRUCTION_SIZE	  : integer;
		SIGN_EXTENSION_SIZE : integer);
	 port (
		clk				: in	std_logic;
		rs1_data			: in	std_logic_vector(REGISTER_SIZE-1 downto 0);
		rs2_data			: in	std_logic_vector(REGISTER_SIZE-1 downto 0);
		current_pc		: in	std_logic_vector(REGISTER_SIZE-1 downto 0);
		predicted_pc	: in	std_logic_vector(REGISTER_SIZE-1 downto 0);
		instr				: in	std_logic_vector(INSTRUCTION_SIZE-1 downto 0);
		sign_extension : in	std_logic_vector(SIGN_EXTENSION_SIZE-1 downto 0);
		data_out			: out std_logic_vector(REGISTER_SIZE-1 downto 0);
		data_out_en		: out std_logic;
		new_pc			: out std_logic_vector(REGISTER_SIZE-1 downto 0);	--next pc
		bad_predict		: out std_logic
		);
  end component branch_unit;

  component load_store_unit is
	 generic (
		REGISTER_SIZE		  : integer;
		SIGN_EXTENSION_SIZE : integer;
		INSTRUCTION_SIZE	  : integer;
		MEMORY_SIZE_BYTES	  : integer);
	 port (
		clk				: in	std_logic;
		valid				: in	std_logic;
		rs1_data			: in	std_logic_vector(REGISTER_SIZE-1 downto 0);
		rs2_data			: in	std_logic_vector(REGISTER_SIZE-1 downto 0);
		instruction		: in	std_logic_vector(INSTRUCTION_SIZE-1 downto 0);
		sign_extension : in	std_logic_vector(SIGN_EXTENSION_SIZE-1 downto 0);
		data_out			: out std_logic_vector(REGISTER_SIZE-1 downto 0);
		data_enable		: out std_logic
		);
  end component load_store_unit;

  signal rs1_data_fwd : std_logic_vector(REGISTER_SIZE-1 downto 0);
  signal rs2_data_fwd : std_logic_vector(REGISTER_SIZE-1 downto 0);

  constant ZERO : std_logic_vector(REGISTER_NAME_SIZE-1 downto 0) := (others => '0');
begin

  --use the previous clock's writeback data when appropriate

  rs1_data_fwd <= wb_data when wb_sel = rs1 and wb_en = '1'and wb_sel /= ZERO else rs1_data;
  rs2_data_fwd <= wb_data when wb_sel = rs2 and wb_en = '1'and wb_sel /= ZERO else rs2_data;

  alu : component arithmetic_unit
	 generic map (
		INSTRUCTION_SIZE	  => INSTRUCTION_SIZE,
		REGISTER_SIZE		  => REGISTER_SIZE,
		SIGN_EXTENSION_SIZE => SIGN_EXTENSION_SIZE)
	 port map (
		clk				=> clk,
		rs1_data			=> rs1_data_fwd,
		rs2_data			=> rs2_data_fwd,
		instruction		=> instruction,
		sign_extension => sign_extension,
		data_out			=> alu_data_out,
		data_enable		=> alu_data_en);


  branch : component branch_unit
	 generic map (
		REGISTER_SIZE		  => REGISTER_SIZE,
		INSTRUCTION_SIZE	  => INSTRUCTION_SIZE,
		SIGN_EXTENSION_SIZE => SIGN_EXTENSION_SIZE)
	 port map(
		clk				=> clk,
		rs1_data			=> rs1_data_fwd,
		rs2_data			=> rs2_data_fwd,
		current_pc		=> pc_current,
		predicted_pc	=> pc_next,
		instr				=> instruction,
		sign_extension => sign_extension,
		data_out			=> br_data_out,
		data_out_en		=> br_data_en,
		new_pc			=> new_pc,
		bad_predict		=> bad_predict);

  ls_unit : component load_store_unit
	 generic map(
		REGISTER_SIZE		  => REGISTER_SIZE,
		SIGN_EXTENSION_SIZE => SIGN_EXTENSION_SIZE,
		INSTRUCTION_SIZE	  => INSTRUCTION_SIZE,
		MEMORY_SIZE_BYTES	  => 1024)
	 port map(
		clk				=> clk,
		valid				=> '1',
		rs1_data			=> rs1_data_fwd,
		rs2_data			=> rs2_data_fwd,
		instruction		=> instruction,
		sign_extension => sign_extension,
		data_out			=> ld_data_out,
		data_enable		=> ld_data_en);


  --the above components have output latches,
  --find out which is the actual output
  writeback_1hot(2) <= alu_data_en;
  writeback_1hot(1) <= br_data_en;
  writeback_1hot(0) <= ld_data_en;

  with writeback_1hot select
	 wb_data <=
	 alu_data_out	  when "100",
	 br_data_out	  when "010",
	 ld_data_out	  when "001",
	 (others => 'X') when others;

  wb_en				<= alu_data_en or br_data_en or ld_data_en;
  predict_corr_en <= bad_predict;
  predict_corr		<= new_pc;

  --wb_sel needs to be latched as well
  wb_sel_proc : process(clk)
  begin
	 if rising_edge(clk) then
		wb_sel <= rd;
	 end if;
  end process;


  end architecture;
