../../wishbone/wb_ram.vhd