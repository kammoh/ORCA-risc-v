../../wishbone/bram.vhd